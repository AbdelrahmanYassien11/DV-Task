//==============================================================================
// File Name   : uart_base_test.sv
// Author      : Abdelrahman Yassien
// Email       : Abdelrahman.Yassien11@gmail.com
// Created On  : 2026-02-03
//
// Description :
//   Base test class for UART verification. Provides common configuration,
//   environment creation, and utility methods for all derived UART tests.
//
// Revision History:
//   0.1 - Initial version
//
// Notes:
//   - All UART tests must extend from this base test
//   - Contains default configuration and build phase logic
//
// Copyright (c) [2026] [Abdelrahman Mohamed Yassien]. All Rights Reserved.
//==============================================================================
`ifndef UART_BASE_TST
`define UART_BASE_TST
class uart_base_test extends uvm_test;
  
  uart_env env;
  uart_config cfg;
  
  `uvm_component_utils(uart_base_test)
  
  function new(string name = "uart_base_test", uvm_component parent = null);
    super.new(name, parent);
  endfunction
  
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    
    // Create configuration
    cfg = uart_config::type_id::create("cfg");
    cfg.set_baud_rate(115200);
    
    // Set configuration in config_db
    uvm_config_db#(uart_config)::set(this, "*", "cfg", cfg);
    
    // Create environment
    env = uart_env::type_id::create("env", this);
  endfunction
  
  function void end_of_elaboration_phase(uvm_phase phase);
    super.end_of_elaboration_phase(phase);
    uvm_top.print_topology();
  endfunction
  
endclass

`endif