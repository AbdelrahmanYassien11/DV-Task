`define TX_DATA_WIDTH 8
`define START_BITS_WIDTH 1
`define STOP_BITS_WIDTH 1
`define PARITY_BITS_WIDTH 1

`define LITERAL(WIDTH, VALUE) WIDTH``'b``VALUE